/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Arkadiusz Kurnik
 * 
 * Description:
 * calculates score for 7seg display
 */

 `timescale 1 ns / 1 ps

 module ctl_score(

 );

 endmodule